module ei_adder32 (
    input [31:0] a,
    input [31:0] b,
    input cin,          
    output [31:0] sum,
    output cout
);
    wire [32:0] c;
    assign c[0] = cin; 

    genvar i;
    generate
        for(i=0; i<32; i=i+1) begin: ADD_LOOP
            full_adder fa (.a(a[i]), .b(b[i]), .cin(c[i]), .sum(sum[i]), .cout(c[i+1]));
        end
    endgenerate
    assign cout = c[32];
endmodule	